`timescale 1ns / 1ps

module Top_Module(
    input clk,              // 100 MHz Sistem Saati
    input rst,              // Reset Butonu (btnC) - Ekran� temizlemek i�in �art!
    input [3:0] col,        // Keypad S�tunlar� (PMOD'dan gelir)
    output [3:0] row,       // Keypad Sat�rlar� (PMOD'a gider)
    output [6:0] seg,       // 7-Segment Segmentler
    output [3:0] an,        // 7-Segment Anotlar
    output dp               // Nokta
    );

    // --- �� KABLOLAR (Wires) ---
    wire w_slow_clk;        // Clock Divider'dan ��kan yava� saat
    wire [3:0] w_key_data;  // Scanner'dan okunan HAFIZALI tu� verisi

    // 1. Mod�l: Saat B�l�c�
    // Scanner'�n h�z�n� belirler (2.5 Milyon / 20Hz civar� idealdir)
    Clock_Divider Divider_Unit (
        .clk(clk),
        .rst(rst),
        .slow_clk(w_slow_clk)
    );

    // 2. Mod�l: Keypad Taray�c� (Yeni Resetli ve Haf�zal� Versiyon)
    // Debouncer olmad��� i�in do�rudan bu mod�lden ��kan veriyi kullanaca��z.
    Keypad_Scanner Scanner_Unit (
        .clk(w_slow_clk),   // Yava� saat
        .rst(rst),          // YEN�: Haf�zay� silmek i�in reset laz�m
        .col(col),          // Giri�
        .row(row),          // ��k��
        .key_out(w_key_data) // Tu� verisi (Bas�lmad���nda son de�eri korur)
    );

    // 3. Mod�l: Ekran S�r�c�
    // Arada Debouncer YOK. Scanner ��k��� direkt buraya giriyor.
    Seven_Seg_Driver Display_Unit (
        .clk(clk),           // 100 MHz (Kombinasyonel oldu�u i�in fark etmez)
        .in_number(w_key_data), // D�KKAT: Direkt w_key_data ba�land�
        .seg(seg),
        .an(an),
        .dp(dp)
    );

endmodule